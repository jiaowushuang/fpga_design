`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name:    sd_write 
//////////////////////////////////////////////////////////////////////////////////
module sd_write(  
		input SD_clk,
		output reg SD_cs,            //SD卡控制器的使能
		output reg SD_datain,
		input  SD_dataout,
						
		input [31:0] sec,            // 写SD的sec地址(注意这是4G内存);且为图像数据地址
									 // 有可能不会作为输入；而是由自己进行配置一个初始值。
		input [31:0] sec_catalog,    // 目录项地址
		
		input write_req,             // 这里没必要存在；控制写的触发条件是根据写使能和一定的延迟决定；
		                             // 而该延迟是COMS照相机的拍照间隔时间。

		output reg rx_valid,         // 接收SD卡的应答响应信号（SD卡是命令/响应型）
						
		input init,                  

		output reg [3:0] mystate,     //状态机的状态可以省略
		output reg write_o            //写使能信号
						
						
    );
	 
	 
	 
//wire [3:0] mystate_o; //调试用
reg [7:0] rx; //FIFO用于将一位的输入数据转换为8位；
//reg [7:0] write_data; //调试用

reg en;          //使能:接受输入的数据
reg [5:0] aa;    //计数等待8个时钟
reg [21:0] cnt;  //写CRC计数16次或是其他计数

reg [47:0] CMD24={8'h58,8'h00,8'h00,8'h00,8'h00,8'hff};//CMD24的字节序列（初始值）
reg [7:0] Sblock_token=8'hfe; //检验块

//reg [7:0] CMDX; //调试用
reg [7:0] CMDY=8'hff; //CRC
reg [2:0] cnta; //计数等待8个时钟

/////////////////////////////   自己定义的参数 
reg flag=0;                     //作为区分两次写操作：一次是写配置文件；一次是写图像数据文件。
								//设置标志位flag，flag=0写入配置文件；flag=1写入图像数据

reg [11:0] sec_size;            //文件的当前长度

reg [31:0] sec_phy= sec_catalog * 512 ;  
								//这里的意思是将sec扇区地址转换为物理地址，便于以后的目录项配置。
								//配置地址寄存器
								
parameter SEC_LEN=12'd3072;     //一张照片的大小（以扇区作为单位） ：1024 * 768 * 2 /512
								//也就是文件的额定长度
								
reg [15:0] delay_cnt;           //作为图像数据发送的延迟

reg [7:0] config_data_reg_0 = 8'bff;   
reg [7:0] config_data_reg_1 = 8'bff; 
reg [7:0] config_data_reg_2 = 8'bff;  
reg [7:0] config_data_reg_3 = 8'bff; 
reg [7:0] config_data_reg_4 = 8'bff; 
reg [7:0] config_data_reg_5 = 8'bff; 
reg [7:0] config_data_reg_06 = 8'bff; 
reg [7:0] config_data_reg_07 = 8'bff; 
reg [7:0] config_data_reg_08 = 8'bff; 
reg [7:0] config_data_reg_09 = 8'bff; 
reg [7:0] config_data_reg_010 = 8'bff; 
reg [7:0] config_data_reg_011 = 8'bff; 
reg [7:0] config_data_reg_012 = 8'bff; 
reg [7:0] config_data_reg_013 = 8'bff; 
reg [7:0] config_data_reg_014 = 8'bff; 
reg [7:0] config_data_reg_015 = 8'bff; 
reg [7:0] config_data_reg_016 = 8'bff; 
reg [7:0] config_data_reg_017 = 8'bff; 
reg [7:0] config_data_reg_018 = 8'bff; 
reg [7:0] config_data_reg_019 = 8'bff; 
reg [7:0] config_data_reg_020 = 8'b00; 

								//作为配置数据的寄存器 ；保守估计有20字节，那就是160位；

reg [7:0]  n=0;                //作为配置文件的角标；由于需要一位一位的配置（SPI模式）

/////////////////////////////状态机的各个状态

parameter idle=4'd0;
parameter write_cmd=4'd1;
parameter wait_8clk=4'd2;
parameter start_r1=4'b3;
parameter start_taken=4'd4;
parameter writea=4'd5;
parameter write_crc=4'd6;
parameter write_wait=4'd7;
parameter write_done=4'd8;


//SD卡写程序
always @(negedge SD_clk)
if(!init)
	begin
	mystate<=idle;
	CMD24<={8'h58,8'h00,8'h00,8'h00,8'h00,8'hff};
	write_o<=1'b0;
	sec_size<=0;
	end
else
	begin
	case(mystate)
		idle:	
		begin
		SD_cs<=1'b1;
		SD_datain<=1'b1;
		cnt<=22'd0;	
		if((write_o==1'b0) && (delay_cnt==10000)) 
		    begin          //如果有写请求			
			mystate<=write_cmd;
				if(flag==0)CMD24<={8'h58,sec_phy[31:24],sec_phy[23:16],sec_phy[15:8],sec_phy[7:0],8'hff};
				else CMD24<={8'h58,sec[31:24],sec[23:16],sec[15:8],sec[7:0],8'hff};
			Sblock_token<=8'hfe;
			write_o<=1'b0;
			end
		else 
		    begin
			mystate<=idle;
			delay_cnt<=delay_cnt+1'b1;	//延迟一秒，每个一秒写一个图像
			end
		end
		
		write_cmd: 
		begin                             //发送CMD24命令 (单块写)	
		if(CMD24!=48'd0) 
		    begin
			SD_cs<=1'b0;
			SD_datain<=CMD24[47];
			CMD24<={CMD24[46:0],1'b0};    //移位输出	
			end
		else 
		    begin 
			mystate<=start_r1;
			end
		end
		start_r1:
		////////////////////////////FIFO程序 
		always @(posedge SD_clk)
			begin
			rx[0]<=SD_dataout;
			rx[7:1]<=rx[6:0];
			end
		//接收SD卡的应答数据
		always @(posedge SD_clk)
			begin
				if(!SD_dataout&&!en)                 //等待SD_dataout为低,SD_dataout为低,开始接收数据
					begin 
					rx_valid<=1'b0; 
					aa<=1;
					en<=1'b1;
					end      
				else if(en)	
					begin 
						if(aa<7) 
							begin
							aa<=aa+1'b1; 
							rx_valid<=1'b0;
							end
						else 
							begin
							aa<=0;
							en<=1'b0;
							rx_valid<=1'b1;             //等待8个CLK后,rx_valid信号开始有效
							end
					end
				else 
					begin 
					cnta<=7;
					SD_cs<=1'b1;	
					en<=1'b0;
					aa<=0;
					rx_valid<=1'b0;
					SD_datain<=1'b1;
					mystate<=wait_8clk;
					end
			end	    
		wait_8clk: 
		begin                            //写数据之前等待8clock
			if(cnta>0) 
			    begin
				cnta<=cnta-1'b1;
				SD_cs<=1'b1;
				SD_datain<=1'b1;
			    end
		    else 
			    begin
			    SD_cs<=1'b1;
				SD_datain<=1'b1;
				mystate<=start_taken;
				cnta<=7;
			    end
				
		end		
		start_taken: 
		begin                           //发送Start Block Taken ：oxfe
			if(cnta>0) 
			    begin
			    cnta<=cnta-1'b1;
				SD_cs<=1'b0;
				SD_datain<=Sblock_token[cnta];
			    end
			else
     			begin
				SD_cs<=1'b0;
				SD_datain<=Sblock_token[0];
				mystate<=writea;
			    cnta<=7;
			    cnt<=0;
				end
		end
//////////////////////////////////////////写文件过程
		writea: 
		begin
//////////////////////////////////////////第一次写配置文件
		    if(flag==0)
			    begin
			    flag<=1;
				
			//配置文件内容
			        if(cnt<512)	
					    begin		
			                if(cnta>=0)	
								begin
				  		        SD_cs<=1'b0;
									if(sec_phy)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_0[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_0[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_0[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_0[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_0[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_0[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_0[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_0[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
							        end
					                else if(sec_phy+1)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_1[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_1[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_1[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_1[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_1[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_1[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_1[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_1[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
						            else if(sec_phy+2)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_2[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_2[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_2[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_2[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_2[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_2[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_2[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_2[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+3)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_3[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_3[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_3[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_3[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_3[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_3[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_3[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_3[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+4)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_4[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_4[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_4[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_4[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_4[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_4[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_4[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_4[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+5)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_5[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_5[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_5[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_5[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_5[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_5[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_5[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_5[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+6)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_06[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_06[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_06[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_06[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_06[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_06[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_06[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_06[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+7)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_07[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_07[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_07[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_07[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_07[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_07[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_07[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_07[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+8)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_08[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_08[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_08[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_08[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_08[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_08[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_08[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_08[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+9)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_09[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_09[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_09[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_09[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_09[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_09[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_09[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_09[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+10)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_010[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_010[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_010[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_010[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_010[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_010[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_010[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_010[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+11)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_011[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_011[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_011[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_011[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_011[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_011[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_011[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_011[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+12)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_012[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_012[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_012[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_012[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_012[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_012[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_012[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_012[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+13)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_013[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_013[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_013[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_013[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_013[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_013[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_013[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_013[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+14)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_014[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_014[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_014[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_014[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_014[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_014[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_014[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_014[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+15)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_015[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_015[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_015[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_015[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_015[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_015[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_015[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_015[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+16)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_016[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_016[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_016[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_016[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_016[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_016[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_016[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_016[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+17)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_017[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_017[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_017[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_017[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_017[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_017[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_017[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_017[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else if(sec_phy+18)
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_018[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_018[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_018[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_018[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_018[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_018[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_018[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_018[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
									else 
									begin
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_019[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_019[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_019[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_019[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_019[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_019[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_019[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_019[7];
						                cnta<=cnta-1'b1;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
						            end
				                end
							else
								begin
									SD_cs<=1'b0;
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_020[0];
						                //cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_020[1];
						                //cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_020[2];
						                //cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_020[3];
						               // cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_020[4];
						                //cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_020[5];
						                //cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_020[6];
						                //cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_020[7];
						                cnta<=7;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
								end
						end
			        else 
						begin              //last byte
						if(cnta>=0)	
							    begin
									SD_cs<=1'b0;
							            case(n)
							            1'b0:
										begin
								        SD_datain<=config_data_reg_020[0];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b1:
										begin
								        SD_datain<=config_data_reg_020[1];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
							            1'b2:
										begin
								        SD_datain<=config_data_reg_020[2];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b3:
										begin
								        SD_datain<=config_data_reg_020[3];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b4:
										begin
								        SD_datain<=config_data_reg_020[4];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b5:
										begin
								        SD_datain<=config_data_reg_020[5];
						                cnta<=cnta-1'b1;
								        n<=n+1;
							            end
										1'b6:
										begin
										SD_datain<=config_data_reg_020[6];
						                cnta<=cnta-1'b1;
								        n<=n+1;
										end
										1'b7:
										begin
										SD_datain<=config_data_reg_020[7];
						                cnta<=cnta-1'b1;
								        n<=0;
										cnt<=cnt+1;
							            default:n<=0;
							            endcase
									sec_phy<=sec_phy+1;
								end
						else 
							begin
							n<=0;
							cnt<=0;
							end	
						end	
					end
				end 
///////////////////////////////////第二次写图像数据				
			else 
				begin             //写512个bytes
				//xxxxxx需要SD_dataout与COMS摄像头的数据线相连；这样需要一个使能信号和COMS信号；这里可以在例化时书写
					if(cnt<512)	
						begin		
							if(cnta>0)	
								begin
								SD_cs<=1'b0;
								SD_datain<=SD_dataout[cnta];
								cnta<=cnta-1'b1;
								end
							else
								begin
								SD_cs<=1'b0;
								SD_datain<=SD_dataout[0];
								cnta<=7;
								cnt<=cnt+1'b1;
								end
						end
					else 
						begin              //last byte
							if(cnta>0)
								begin
								SD_datain<=SD_dataout[cnta];
								cnta<=cnta-1'b1;
								end
							else 
								begin
								SD_datain<=SD_dataout[cnta];
								cnta<=7;
								cnt<=0;
								mystate<=write_crc;						
								end
						end
				end
		end

///////////////////////////////////////////////////////////////////
		write_crc: 
		begin               //写crc:0xff
				if(cnt<16) 
				    begin
					SD_cs<=1'b0;
					SD_datain<=1'b1;
					cnt<=cnt+1'b1;
				    end
				else 
				    begin
				    if(rx_valid)         //等待Data Response Token
						mystate<=write_wait;
					else
					    mystate<=write_crc;					 
				    end
		end
		write_wait: 
		begin               //等待数据写入完成
		    if(rx==8'hxx)   //改为正确的RX值或是有值即可
			    begin
					mystate<=write_done;	 
				end
			else 
			    begin 
					mystate<=write_wait;
				end
		end
		write_done:
		begin
			if(cnt<22'd15)
     			begin      //等待15个clock
				SD_cs<=1'b1;
				SD_datain<=1'b1;
				cnt<=cnt+1'b1;
			    end
			else
     			begin  
				cnt<=0;
					if (sec_size<SEC_LEN) 
					    begin                           //如果整幅图像还未写完 
 					    write_o<=1'b0;
                        sec <= sec + 1;                 //加1，即为512字节
						sec_size <= sec_size +1;
						mystate<=idle;
					    end	 
					else	
					    begin	 
					    write_o<=1'b1;
						mystate<=idle;
					    end	 

				end					
		end		
		default:mystate<=idle;
		endcase		
	end					
endmodule
